magic
tech sky130A
magscale 1 2
timestamp 1729047055
<< error_p >>
rect -136 -1229 -78 -1223
rect 655 -1229 713 -1223
rect 1446 -1229 1504 -1223
rect -136 -1263 -124 -1229
rect 655 -1263 667 -1229
rect 1446 -1263 1458 -1229
rect -136 -1269 -78 -1263
rect 655 -1269 713 -1263
rect 1446 -1269 1504 -1263
rect -180 -1362 -168 -1350
rect -134 -1362 -80 -1350
rect -46 -1362 -34 -1350
rect 34 -1361 68 -1343
rect 34 -1362 104 -1361
rect -205 -1384 -180 -1362
rect -168 -1370 -9 -1362
rect -205 -1388 -168 -1384
rect -134 -1388 -9 -1370
rect -205 -1396 -9 -1388
rect 33 -1397 104 -1362
rect -177 -1448 -168 -1414
rect -143 -1426 -122 -1417
rect -92 -1426 -77 -1417
rect -165 -1447 -122 -1426
rect -165 -1448 -121 -1447
rect -93 -1448 -55 -1426
rect -46 -1448 -43 -1414
rect 51 -1431 122 -1397
rect -165 -1454 -132 -1448
rect -123 -1449 -122 -1448
rect -93 -1454 -34 -1448
rect -165 -1482 -34 -1454
rect -180 -1489 -34 -1482
rect -193 -1501 -27 -1489
rect -168 -1505 -45 -1501
rect -160 -1515 -45 -1505
rect -143 -1523 -45 -1515
rect -143 -1532 -40 -1523
rect -171 -1536 -40 -1532
rect 51 -1533 121 -1431
rect 279 -1483 295 -1326
rect 470 -1456 473 -1361
rect 611 -1362 623 -1350
rect 657 -1362 711 -1350
rect 745 -1362 757 -1350
rect 825 -1361 859 -1343
rect 825 -1362 895 -1361
rect 586 -1384 611 -1362
rect 623 -1370 782 -1362
rect 586 -1388 623 -1384
rect 657 -1388 782 -1370
rect 586 -1396 782 -1388
rect 824 -1397 895 -1362
rect 614 -1438 623 -1414
rect 648 -1426 669 -1417
rect 699 -1426 714 -1417
rect 611 -1448 623 -1438
rect 626 -1447 669 -1426
rect 626 -1448 670 -1447
rect 698 -1448 736 -1426
rect 745 -1448 748 -1414
rect 842 -1431 913 -1397
rect 611 -1454 659 -1448
rect 668 -1449 669 -1448
rect 698 -1454 757 -1448
rect 611 -1456 757 -1454
rect 470 -1489 757 -1456
rect 235 -1490 289 -1489
rect 235 -1492 295 -1490
rect 235 -1493 441 -1492
rect 233 -1499 441 -1493
rect 197 -1511 277 -1499
rect 279 -1511 441 -1499
rect 197 -1526 441 -1511
rect 197 -1533 283 -1526
rect -190 -1598 -183 -1536
rect -171 -1537 -137 -1536
rect -95 -1537 -90 -1536
rect -83 -1537 -49 -1536
rect -171 -1539 -126 -1537
rect -95 -1539 -49 -1537
rect -143 -1548 -126 -1539
rect -187 -1616 -183 -1598
rect -162 -1588 -126 -1548
rect -124 -1548 -60 -1539
rect -124 -1573 -52 -1548
rect -95 -1574 -94 -1573
rect -91 -1574 -90 -1573
rect -162 -1589 -125 -1588
rect -95 -1589 -94 -1588
rect -83 -1589 -52 -1573
rect -162 -1590 -124 -1589
rect -96 -1590 -52 -1589
rect -162 -1607 -125 -1590
rect -171 -1611 -125 -1607
rect -171 -1616 -149 -1611
rect -187 -1639 -149 -1616
rect -140 -1620 -125 -1611
rect -95 -1607 -52 -1590
rect -37 -1598 -24 -1536
rect 51 -1539 291 -1533
rect 51 -1549 283 -1539
rect 295 -1549 441 -1526
rect 470 -1501 764 -1489
rect 470 -1505 746 -1501
rect 470 -1532 627 -1505
rect 631 -1515 746 -1505
rect 648 -1523 746 -1515
rect 648 -1532 751 -1523
rect 470 -1536 751 -1532
rect 842 -1533 912 -1431
rect 1070 -1483 1086 -1326
rect 1261 -1456 1264 -1361
rect 1402 -1362 1414 -1350
rect 1448 -1362 1502 -1350
rect 1536 -1362 1548 -1350
rect 1616 -1361 1650 -1343
rect 1616 -1362 1686 -1361
rect 1377 -1384 1402 -1362
rect 1414 -1370 1573 -1362
rect 1377 -1388 1414 -1384
rect 1448 -1388 1573 -1370
rect 1377 -1396 1573 -1388
rect 1615 -1397 1686 -1362
rect 1405 -1438 1414 -1414
rect 1439 -1426 1460 -1417
rect 1490 -1426 1505 -1417
rect 1402 -1448 1414 -1438
rect 1417 -1447 1460 -1426
rect 1417 -1448 1461 -1447
rect 1489 -1448 1527 -1426
rect 1536 -1448 1539 -1414
rect 1633 -1431 1704 -1397
rect 1402 -1454 1450 -1448
rect 1459 -1449 1460 -1448
rect 1489 -1454 1548 -1448
rect 1402 -1456 1548 -1454
rect 1261 -1489 1548 -1456
rect 1026 -1490 1080 -1489
rect 1026 -1492 1086 -1490
rect 1026 -1493 1232 -1492
rect 1024 -1499 1232 -1493
rect 988 -1511 1068 -1499
rect 1070 -1511 1232 -1499
rect 988 -1526 1232 -1511
rect 988 -1533 1074 -1526
rect 470 -1537 654 -1536
rect 696 -1537 701 -1536
rect 708 -1537 742 -1536
rect 470 -1539 665 -1537
rect 696 -1539 742 -1537
rect 470 -1548 645 -1539
rect 648 -1548 665 -1539
rect 51 -1576 297 -1549
rect 51 -1580 309 -1576
rect -95 -1611 -49 -1607
rect -95 -1620 -74 -1611
rect -71 -1616 -49 -1611
rect -37 -1616 -33 -1598
rect -183 -1675 -149 -1639
rect -71 -1639 -33 -1616
rect -71 -1641 -37 -1639
rect -61 -1675 -49 -1641
rect -37 -1675 -3 -1641
rect 51 -1675 121 -1580
rect 207 -1605 309 -1580
rect 403 -1588 414 -1567
rect 426 -1588 437 -1567
rect 470 -1588 665 -1548
rect 667 -1548 731 -1539
rect 667 -1573 739 -1548
rect 696 -1574 697 -1573
rect 700 -1574 701 -1573
rect -183 -1700 -158 -1675
rect -62 -1700 -37 -1675
rect -139 -1774 -81 -1768
rect -139 -1808 -127 -1774
rect -139 -1814 -81 -1808
rect 51 -1910 119 -1675
rect 207 -1755 235 -1605
rect 241 -1621 309 -1605
rect 387 -1594 445 -1588
rect 470 -1589 666 -1588
rect 696 -1589 697 -1588
rect 708 -1589 739 -1573
rect 470 -1590 667 -1589
rect 695 -1590 739 -1589
rect 241 -1675 335 -1621
rect 387 -1628 399 -1594
rect 403 -1628 437 -1594
rect 470 -1611 666 -1590
rect 387 -1634 445 -1628
rect 355 -1675 357 -1671
rect 369 -1675 389 -1671
rect 241 -1692 309 -1675
rect 241 -1755 275 -1692
rect 207 -1780 275 -1755
rect 207 -1784 235 -1780
rect 241 -1818 275 -1780
rect 289 -1784 309 -1692
rect 317 -1768 329 -1675
rect 321 -1780 329 -1768
rect 343 -1763 389 -1675
rect 403 -1675 437 -1634
rect 470 -1641 645 -1611
rect 651 -1620 666 -1611
rect 696 -1607 739 -1590
rect 754 -1598 767 -1536
rect 842 -1539 1082 -1533
rect 842 -1549 1074 -1539
rect 1086 -1549 1232 -1526
rect 1261 -1501 1555 -1489
rect 1261 -1505 1537 -1501
rect 1261 -1532 1418 -1505
rect 1422 -1515 1537 -1505
rect 1439 -1523 1537 -1515
rect 1439 -1532 1542 -1523
rect 1261 -1536 1542 -1532
rect 1633 -1533 1703 -1431
rect 1861 -1483 1877 -1326
rect 1817 -1490 1871 -1489
rect 1817 -1492 1877 -1490
rect 1817 -1493 2023 -1492
rect 1815 -1499 2023 -1493
rect 1779 -1511 1859 -1499
rect 1861 -1511 2023 -1499
rect 1779 -1526 2023 -1511
rect 1779 -1533 1865 -1526
rect 1261 -1537 1445 -1536
rect 1487 -1537 1492 -1536
rect 1499 -1537 1533 -1536
rect 1261 -1539 1456 -1537
rect 1487 -1539 1533 -1537
rect 1261 -1548 1436 -1539
rect 1439 -1548 1456 -1539
rect 842 -1576 1088 -1549
rect 842 -1580 1100 -1576
rect 696 -1611 742 -1607
rect 696 -1620 717 -1611
rect 720 -1616 742 -1611
rect 754 -1616 758 -1598
rect 720 -1639 758 -1616
rect 720 -1641 754 -1639
rect 470 -1671 642 -1641
rect 443 -1675 642 -1671
rect 730 -1675 742 -1641
rect 754 -1675 788 -1641
rect 842 -1675 912 -1580
rect 998 -1605 1100 -1580
rect 1194 -1588 1205 -1567
rect 1217 -1588 1228 -1567
rect 1261 -1588 1456 -1548
rect 1458 -1548 1522 -1539
rect 1458 -1573 1530 -1548
rect 1487 -1574 1488 -1573
rect 1491 -1574 1492 -1573
rect 403 -1736 645 -1675
rect 729 -1700 754 -1675
rect 403 -1763 627 -1736
rect 343 -1780 627 -1763
rect 321 -1784 323 -1780
rect 349 -1806 361 -1780
rect 349 -1808 357 -1806
rect 355 -1818 357 -1808
rect 241 -1821 265 -1818
rect 233 -1827 291 -1821
rect 233 -1835 265 -1827
rect 233 -1853 245 -1835
rect 275 -1853 279 -1839
rect 233 -1861 279 -1853
rect 233 -1867 291 -1861
rect 369 -1867 627 -1780
rect 652 -1774 710 -1768
rect 652 -1808 664 -1774
rect 652 -1814 710 -1808
rect 241 -1888 275 -1867
rect 357 -1875 627 -1867
rect 369 -1879 627 -1875
rect 381 -1892 627 -1879
rect 373 -1906 627 -1892
rect 51 -1946 101 -1910
rect 237 -1913 627 -1906
rect 237 -1914 403 -1913
rect 237 -1916 433 -1914
rect 437 -1916 627 -1913
rect 237 -1922 627 -1916
rect 237 -1923 434 -1922
rect 237 -1929 433 -1923
rect 437 -1929 627 -1922
rect 237 -1946 627 -1929
rect 842 -1910 910 -1675
rect 998 -1755 1026 -1605
rect 1032 -1621 1100 -1605
rect 1178 -1594 1236 -1588
rect 1261 -1589 1457 -1588
rect 1487 -1589 1488 -1588
rect 1499 -1589 1530 -1573
rect 1261 -1590 1458 -1589
rect 1486 -1590 1530 -1589
rect 1032 -1675 1126 -1621
rect 1178 -1628 1190 -1594
rect 1194 -1628 1228 -1594
rect 1261 -1611 1457 -1590
rect 1178 -1634 1236 -1628
rect 1146 -1675 1148 -1671
rect 1160 -1675 1180 -1671
rect 1032 -1692 1100 -1675
rect 1032 -1755 1066 -1692
rect 998 -1780 1066 -1755
rect 998 -1784 1026 -1780
rect 1032 -1818 1066 -1780
rect 1080 -1784 1100 -1692
rect 1108 -1768 1120 -1675
rect 1112 -1780 1120 -1768
rect 1134 -1763 1180 -1675
rect 1194 -1675 1228 -1634
rect 1261 -1641 1436 -1611
rect 1442 -1620 1457 -1611
rect 1487 -1607 1530 -1590
rect 1545 -1598 1558 -1536
rect 1633 -1539 1873 -1533
rect 1633 -1549 1865 -1539
rect 1877 -1549 2023 -1526
rect 1633 -1576 1879 -1549
rect 1633 -1580 1891 -1576
rect 1487 -1611 1533 -1607
rect 1487 -1620 1508 -1611
rect 1511 -1616 1533 -1611
rect 1545 -1616 1549 -1598
rect 1511 -1639 1549 -1616
rect 1511 -1641 1545 -1639
rect 1261 -1671 1433 -1641
rect 1234 -1675 1433 -1671
rect 1521 -1675 1533 -1641
rect 1545 -1675 1579 -1641
rect 1633 -1675 1703 -1580
rect 1789 -1605 1891 -1580
rect 1985 -1588 1996 -1567
rect 2008 -1588 2019 -1567
rect 1194 -1736 1436 -1675
rect 1520 -1700 1545 -1675
rect 1194 -1763 1418 -1736
rect 1134 -1780 1418 -1763
rect 1112 -1784 1114 -1780
rect 1140 -1806 1152 -1780
rect 1140 -1808 1148 -1806
rect 1146 -1818 1148 -1808
rect 1032 -1821 1056 -1818
rect 1024 -1827 1082 -1821
rect 1024 -1835 1056 -1827
rect 1024 -1853 1036 -1835
rect 1066 -1853 1070 -1839
rect 1024 -1861 1070 -1853
rect 1024 -1867 1082 -1861
rect 1160 -1867 1418 -1780
rect 1443 -1774 1501 -1768
rect 1443 -1808 1455 -1774
rect 1443 -1814 1501 -1808
rect 1032 -1888 1066 -1867
rect 1148 -1875 1418 -1867
rect 1160 -1879 1418 -1875
rect 1172 -1892 1418 -1879
rect 1164 -1906 1418 -1892
rect 842 -1946 892 -1910
rect 1028 -1913 1418 -1906
rect 1028 -1914 1194 -1913
rect 1028 -1916 1224 -1914
rect 1228 -1916 1418 -1913
rect 1028 -1922 1418 -1916
rect 1028 -1923 1225 -1922
rect 1028 -1929 1224 -1923
rect 1228 -1929 1418 -1922
rect 1028 -1946 1418 -1929
rect 1633 -1910 1701 -1675
rect 1789 -1755 1817 -1605
rect 1823 -1621 1891 -1605
rect 1969 -1594 2027 -1588
rect 1823 -1675 1917 -1621
rect 1969 -1628 1981 -1594
rect 1985 -1628 2019 -1594
rect 1969 -1634 2027 -1628
rect 1937 -1675 1939 -1671
rect 1951 -1675 1971 -1671
rect 1823 -1692 1891 -1675
rect 1823 -1755 1857 -1692
rect 1789 -1780 1857 -1755
rect 1789 -1784 1817 -1780
rect 1823 -1818 1857 -1780
rect 1871 -1784 1891 -1692
rect 1899 -1768 1911 -1675
rect 1903 -1780 1911 -1768
rect 1925 -1763 1971 -1675
rect 1985 -1675 2019 -1634
rect 2025 -1675 2053 -1671
rect 1985 -1763 2053 -1675
rect 1925 -1780 2053 -1763
rect 1903 -1784 1905 -1780
rect 1931 -1806 1943 -1780
rect 1931 -1808 1939 -1806
rect 1937 -1818 1939 -1808
rect 1823 -1821 1847 -1818
rect 1815 -1827 1873 -1821
rect 1951 -1825 2053 -1780
rect 1815 -1835 1847 -1827
rect 1815 -1853 1827 -1835
rect 1857 -1853 1861 -1839
rect 1815 -1861 1861 -1853
rect 1815 -1867 1873 -1861
rect 1951 -1867 2063 -1825
rect 1823 -1888 1857 -1867
rect 1939 -1875 2063 -1867
rect 1951 -1879 2185 -1875
rect 1963 -1892 2185 -1879
rect 1955 -1906 2185 -1892
rect 1633 -1946 1683 -1910
rect 1819 -1913 2185 -1906
rect 1819 -1914 1985 -1913
rect 1819 -1916 2015 -1914
rect 2019 -1916 2185 -1913
rect 1819 -1922 2185 -1916
rect 1819 -1923 2016 -1922
rect 1819 -1929 2015 -1923
rect 2019 -1929 2065 -1922
rect 237 -1962 483 -1946
rect 237 -1963 391 -1962
rect 437 -1963 483 -1962
rect 383 -1972 483 -1963
rect 383 -2006 449 -1972
rect 842 -1999 881 -1946
rect 1028 -1962 1274 -1946
rect 1028 -1963 1182 -1962
rect 1228 -1963 1274 -1962
rect 1174 -1972 1274 -1963
rect 1174 -2006 1240 -1972
rect 1633 -1999 1672 -1946
rect 1819 -1962 2065 -1929
rect 1819 -1963 1973 -1962
rect 2019 -1963 2065 -1962
rect 1965 -1972 2065 -1963
rect 1965 -2006 2031 -1972
rect 383 -2129 399 -2006
rect 1174 -2129 1190 -2006
rect 1965 -2129 1981 -2006
use ring_osilator  x1
timestamp 1729047055
transform 1 0 0 0 1 -833
box -321 -1296 2209 2550
<< end >>
