magic
tech sky130A
magscale 1 2
timestamp 1729327972
<< nwell >>
rect -1456 2322 797 3540
<< viali >>
rect -628 3470 -594 3504
rect -9 3470 343 3504
<< metal1 >>
rect -695 3504 388 3529
rect -695 3470 -628 3504
rect -594 3470 -9 3504
rect 343 3470 388 3504
rect -695 3456 388 3470
rect 521 2960 573 2966
rect -474 2915 44 2949
rect -643 2779 -637 2831
rect -585 2822 -579 2831
rect -474 2822 -440 2915
rect 521 2902 573 2908
rect -585 2788 -440 2822
rect -585 2779 -579 2788
rect -351 2299 -345 2359
rect -285 2299 -279 2359
rect -722 2169 -477 2217
rect -332 2173 -298 2299
rect -541 602 -477 2169
rect -110 1213 240 1359
rect -207 1038 -201 1098
rect -141 1038 -135 1098
rect -547 538 -541 602
rect -477 538 -471 602
rect 111 -195 117 -143
rect 169 -195 175 -143
<< via1 >>
rect -637 2779 -585 2831
rect 521 2908 573 2960
rect -345 2299 -285 2359
rect -201 1038 -141 1098
rect -541 538 -477 602
rect 117 -195 169 -143
<< metal2 >>
rect -234 2960 -178 2969
rect 515 2951 521 2960
rect 372 2917 521 2951
rect 515 2908 521 2917
rect 573 2908 579 2960
rect -234 2895 -178 2904
rect -637 2831 -585 2837
rect -637 2773 -585 2779
rect 857 2466 913 2475
rect 234 2421 857 2455
rect 857 2401 913 2410
rect -345 2359 -285 2365
rect -352 2301 -345 2357
rect -285 2301 -278 2357
rect -345 2293 -285 2299
rect -998 2078 -989 2138
rect -929 2078 -920 2138
rect -534 2136 -474 2138
rect -541 2080 -532 2136
rect -476 2080 -467 2136
rect -534 1303 -474 2080
rect 606 1769 615 1829
rect 675 1769 684 1829
rect -534 1243 -141 1303
rect -201 1098 -141 1243
rect -201 1032 -141 1038
rect -541 602 -477 608
rect -541 532 -477 538
rect 117 -143 169 45
rect 117 -201 169 -195
<< via2 >>
rect -234 2904 -178 2960
rect 857 2410 913 2466
rect -343 2301 -287 2357
rect -989 2078 -929 2138
rect -532 2080 -476 2136
rect 615 1769 675 1829
rect -537 542 -481 598
<< metal3 >>
rect -239 2962 -173 2965
rect -239 2960 23 2962
rect -239 2904 -234 2960
rect -178 2904 23 2960
rect -239 2902 23 2904
rect -239 2899 -173 2902
rect -348 2359 -282 2362
rect 155 2359 215 2468
rect 852 2466 918 2471
rect 852 2410 857 2466
rect 913 2410 918 2466
rect 852 2405 918 2410
rect -348 2357 215 2359
rect -348 2301 -343 2357
rect -287 2301 215 2357
rect -348 2299 215 2301
rect -348 2296 -282 2299
rect -994 2138 -924 2143
rect -537 2138 -471 2141
rect -994 2078 -989 2138
rect -929 2136 -471 2138
rect -929 2080 -532 2136
rect -476 2080 -471 2136
rect -929 2078 -471 2080
rect -994 2073 -924 2078
rect -537 2075 -471 2078
rect 610 1829 680 1834
rect 855 1829 915 2405
rect 610 1769 615 1829
rect 675 1769 915 1829
rect 610 1764 680 1769
rect -542 602 -476 603
rect -542 598 -81 602
rect -542 542 -537 598
rect -481 542 -81 598
rect -542 538 -81 542
rect -542 537 -476 538
use NMOS34  NMOS34_0 ~/mag/NMOS34
timestamp 1729215808
transform 1 0 -140 0 1 -53
box -292 -71 973 1317
use NMOS89  NMOS89_0 ~/mag/NMOS89
timestamp 1729222480
transform 1 0 -256 0 1 1377
box -176 -71 1106 917
use PMOS67  PMOS67_0 ~/mag/PMOS67
timestamp 1729239979
transform 1 0 -190 0 1 1495
box -267 827 987 2045
use PMOS125  PMOS125_0 ~/mag/PMOS125
timestamp 1729186466
transform 1 0 -1251 0 1 817
box -205 -139 793 2723
<< labels >>
flabel metal1 -288 3487 -288 3487 0 FreeSans 800 0 0 0 VDD
port 1 nsew
flabel metal1 50 1287 51 1287 0 FreeSans 800 0 0 0 GND
port 2 nsew
flabel metal3 883 2243 883 2243 0 FreeSans 800 0 0 0 OUT
port 3 nsew
flabel via1 145 -167 145 -167 0 FreeSans 800 0 0 0 RS
port 6 nsew
flabel via2 -208 2934 -206 2935 0 FreeSans 800 0 0 0 VIP
port 8 nsew
flabel via1 550 2935 550 2935 0 FreeSans 800 0 0 0 VIN
port 10 nsew
<< end >>
