magic
tech sky130A
magscale 1 2
timestamp 1729186466
<< nwell >>
rect -205 2353 793 2723
rect -205 2296 127 2353
rect 199 2296 793 2353
rect -205 1677 793 2296
rect -205 1666 520 1677
rect -205 1664 233 1666
rect -205 1588 -78 1664
rect 71 1662 233 1664
rect 71 1605 124 1662
rect 196 1605 233 1662
rect 71 1588 233 1605
rect -205 1586 233 1588
rect 336 1663 520 1666
rect 336 1606 387 1663
rect 459 1606 520 1663
rect 336 1593 520 1606
rect 696 1593 793 1677
rect 336 1586 793 1593
rect -205 967 793 1586
rect -205 959 272 967
rect -205 958 124 959
rect -205 895 -70 958
rect 53 902 124 958
rect 196 910 272 959
rect 344 965 518 967
rect 344 910 388 965
rect 196 908 388 910
rect 460 908 518 965
rect 196 902 518 908
rect 53 901 518 902
rect 669 901 793 967
rect 53 895 793 901
rect -205 300 793 895
rect -205 180 -73 300
rect 684 180 793 300
rect -205 -139 793 180
<< nsubdiff >>
rect -169 2653 -109 2687
rect 697 2653 757 2687
rect -169 2627 -135 2653
rect 723 2627 757 2653
rect -169 -69 -135 -43
rect 723 -69 757 -43
rect -169 -103 -109 -69
rect 697 -103 757 -69
<< nsubdiffcont >>
rect -109 2653 697 2687
rect -169 -43 -135 2627
rect 723 -43 757 2627
rect -109 -103 697 -69
<< poly >>
rect -85 2615 7 2631
rect -85 2581 -69 2615
rect -35 2581 7 2615
rect -85 2565 7 2581
rect -23 2533 7 2565
rect 581 2615 673 2631
rect 581 2581 623 2615
rect 657 2581 673 2615
rect 581 2565 673 2581
rect 581 2533 611 2565
rect -85 1921 7 1937
rect 65 1936 265 2036
rect -85 1887 -69 1921
rect -35 1887 7 1921
rect -85 1871 7 1887
rect -23 1839 7 1871
rect 581 1921 673 1937
rect 581 1887 623 1921
rect 657 1887 673 1921
rect 581 1871 673 1887
rect 581 1839 611 1871
rect 65 1242 523 1342
rect -23 713 7 745
rect -85 697 7 713
rect -85 663 -69 697
rect -35 663 7 697
rect -85 647 7 663
rect 581 713 611 745
rect 581 697 673 713
rect 581 663 623 697
rect 657 663 673 697
rect 323 548 523 648
rect 581 647 673 663
rect -23 19 7 51
rect -85 3 7 19
rect -85 -31 -69 3
rect -35 -31 7 3
rect -85 -47 7 -31
rect 581 19 611 51
rect 581 3 673 19
rect 581 -31 623 3
rect 657 -31 673 3
rect 581 -47 673 -31
<< polycont >>
rect -69 2581 -35 2615
rect 623 2581 657 2615
rect -69 1887 -35 1921
rect 623 1887 657 1921
rect -69 663 -35 697
rect 623 663 657 697
rect -69 -31 -35 3
rect 623 -31 657 3
<< locali >>
rect -169 2653 -109 2687
rect 697 2653 757 2687
rect -169 2627 -135 2653
rect 723 2627 757 2653
rect -85 2581 -69 2615
rect -35 2581 -19 2615
rect 607 2581 623 2615
rect 657 2581 673 2615
rect -69 2533 -35 2581
rect 623 2521 657 2581
rect -85 1887 -69 1921
rect -35 1887 -19 1921
rect 607 1887 623 1921
rect 657 1887 673 1921
rect -69 1839 -35 1887
rect 623 1839 657 1887
rect -69 697 -35 745
rect 623 697 657 745
rect -85 663 -69 697
rect -35 663 -19 697
rect 607 663 623 697
rect 657 663 673 697
rect -69 3 -35 51
rect 623 3 657 51
rect -85 -31 -69 3
rect -35 -31 -19 3
rect 607 -31 623 3
rect 657 -31 673 3
rect -169 -69 -135 -43
rect 723 -69 757 -43
rect -169 -103 -109 -69
rect 697 -103 757 -69
<< viali >>
rect 623 2653 657 2687
rect -69 2581 -35 2615
rect 623 2581 657 2615
rect -69 1887 -35 1921
rect 623 1887 657 1921
rect -69 663 -35 697
rect 623 663 657 697
rect -69 -31 -35 3
rect 623 -31 657 3
rect -69 -103 -35 -69
<< metal1 >>
rect 611 2687 669 2693
rect 611 2653 623 2687
rect 657 2653 669 2687
rect -81 2615 -23 2621
rect -81 2581 -69 2615
rect -35 2581 -23 2615
rect -81 2575 -23 2581
rect 611 2615 669 2653
rect 611 2581 623 2615
rect 657 2581 669 2615
rect 611 2575 669 2581
rect -75 2533 -29 2575
rect -88 2133 -78 2533
rect -26 2133 59 2533
rect 271 2092 317 2537
rect 617 2533 663 2575
rect 529 2133 663 2533
rect 529 2092 575 2133
rect 271 2086 382 2092
rect 271 2052 383 2086
rect 271 2046 382 2052
rect 471 2046 575 2092
rect -81 1921 -23 1927
rect -81 1887 -69 1921
rect -35 1887 -23 1921
rect -81 1881 -23 1887
rect -75 1839 -29 1881
rect -75 1439 10 1839
rect 62 1439 72 1839
rect 13 1186 132 1232
rect 13 1145 59 1186
rect -75 745 59 1145
rect -75 703 -29 745
rect -81 697 -23 703
rect -81 663 -69 697
rect -35 663 -23 697
rect -81 657 -23 663
rect 271 538 317 2046
rect 611 1921 669 1927
rect 611 1887 623 1921
rect 657 1887 669 1921
rect 611 1881 669 1887
rect 617 1839 663 1881
rect 529 1439 663 1839
rect 529 1398 575 1439
rect 472 1352 575 1398
rect 516 745 526 1145
rect 578 745 663 1145
rect 617 703 663 745
rect 611 697 669 703
rect 611 663 623 697
rect 657 663 669 697
rect 611 657 669 663
rect 13 492 128 538
rect 211 492 317 538
rect 13 451 59 492
rect -75 51 59 451
rect -75 9 -29 51
rect 271 47 317 492
rect 529 51 614 451
rect 666 51 676 451
rect 617 9 663 51
rect -81 3 -23 9
rect -81 -31 -69 3
rect -35 -31 -23 3
rect -81 -69 -23 -31
rect 611 3 669 9
rect 611 -31 623 3
rect 657 -31 669 3
rect 611 -37 669 -31
rect -81 -103 -69 -69
rect -35 -103 -23 -69
rect -81 -109 -23 -103
<< via1 >>
rect -78 2133 -26 2533
rect 10 1439 62 1839
rect 526 745 578 1145
rect 614 51 666 451
<< metal2 >>
rect -78 2533 -26 2543
rect -78 2123 -26 2133
rect -75 2017 -29 2123
rect -91 1957 -82 2017
rect -22 1957 -13 2017
rect 612 2015 668 2024
rect -75 636 -29 1957
rect 612 1950 668 1959
rect 10 1839 62 1849
rect 10 1317 62 1439
rect 10 1265 578 1317
rect 526 1145 578 1265
rect 526 735 578 745
rect -80 627 -24 636
rect 617 629 663 1950
rect -80 562 -24 571
rect 601 569 610 629
rect 670 569 679 629
rect 617 461 663 569
rect 614 451 666 461
rect 614 41 666 51
<< via2 >>
rect -82 1957 -22 2017
rect 612 1959 668 2015
rect -80 571 -24 627
rect 610 569 670 629
<< metal3 >>
rect -87 2017 -17 2022
rect 607 2017 673 2020
rect -87 1957 -82 2017
rect -22 2015 673 2017
rect -22 1959 612 2015
rect 668 1959 673 2015
rect -22 1957 673 1959
rect -87 1952 -17 1957
rect 607 1954 673 1957
rect -85 629 -19 632
rect 605 629 675 634
rect -85 627 610 629
rect -85 571 -80 627
rect -24 571 610 627
rect -85 569 610 571
rect 670 569 675 629
rect -85 566 -19 569
rect 605 564 675 569
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_0
timestamp 1729132732
transform 1 0 596 0 1 945
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_1
timestamp 1729132732
transform 1 0 596 0 1 2333
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_2
timestamp 1729132732
transform 1 0 -8 0 1 2333
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_3
timestamp 1729132732
transform 1 0 -8 0 1 945
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_4
timestamp 1729132732
transform 1 0 -8 0 1 251
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_5
timestamp 1729132732
transform 1 0 596 0 1 251
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_6
timestamp 1729132732
transform 1 0 596 0 1 1639
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_7
timestamp 1729132732
transform 1 0 -8 0 1 1639
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_0
timestamp 1729185329
transform 1 0 294 0 1 2333
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_1
timestamp 1729185329
transform 1 0 294 0 1 1639
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_2
timestamp 1729185329
transform 1 0 294 0 1 945
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_3
timestamp 1729185329
transform 1 0 294 0 1 251
box -323 -300 323 300
<< labels >>
flabel metal1 640 2635 640 2635 0 FreeSans 160 0 0 0 VDD
port 1 nsew
flabel metal2 641 1290 641 1290 0 FreeSans 160 0 0 0 D5
port 2 nsew
flabel metal1 552 1378 552 1378 0 FreeSans 160 0 0 0 D2
port 3 nsew
flabel metal2 36 1293 36 1293 0 FreeSans 160 0 0 0 D1
port 4 nsew
<< end >>
