magic
tech sky130A
magscale 1 2
timestamp 1729215808
<< psubdiff >>
rect -292 1277 -218 1311
rect 902 1277 973 1311
rect -292 1248 -258 1277
rect 939 1248 973 1277
rect -292 -31 -258 -6
rect 939 -31 973 -6
rect -292 -65 -218 -31
rect 902 -65 973 -31
<< psubdiffcont >>
rect -218 1277 902 1311
rect -292 -6 -258 1248
rect 939 -6 973 1248
rect -218 -65 902 -31
<< poly >>
rect -208 1230 -116 1246
rect -208 1196 -192 1230
rect -158 1196 -116 1230
rect -208 1180 -116 1196
rect -146 1158 -116 1180
rect 797 1230 889 1246
rect 797 1196 839 1230
rect 873 1196 889 1230
rect 797 1180 889 1196
rect 797 1158 827 1180
rect 54 576 626 670
rect -146 66 -116 88
rect -208 50 -116 66
rect -208 16 -192 50
rect -158 16 -116 50
rect -208 0 -116 16
rect 796 66 826 88
rect 796 50 888 66
rect 796 16 838 50
rect 872 16 888 50
rect 796 0 888 16
<< polycont >>
rect -192 1196 -158 1230
rect 839 1196 873 1230
rect -192 16 -158 50
rect 838 16 872 50
<< locali >>
rect -292 1277 -218 1311
rect 902 1277 973 1311
rect -292 1248 -258 1277
rect 939 1248 973 1277
rect -208 1196 -192 1230
rect -158 1196 -142 1230
rect 823 1196 839 1230
rect 873 1196 889 1230
rect -192 1158 -158 1196
rect 839 1158 873 1196
rect -192 50 -158 88
rect 838 50 872 88
rect -208 16 -192 50
rect -158 16 -142 50
rect 822 16 838 50
rect 872 16 888 50
rect -292 -31 -258 -6
rect 939 -31 973 -6
rect -292 -65 -218 -31
rect 902 -65 973 -31
<< viali >>
rect 266 1277 300 1311
rect -192 1196 -158 1230
rect 839 1196 873 1230
rect -192 16 -158 50
rect 838 16 872 50
rect 380 -65 414 -31
<< metal1 >>
rect 254 1311 312 1317
rect 254 1277 266 1311
rect 300 1277 312 1311
rect 254 1271 312 1277
rect -204 1230 -146 1236
rect -204 1196 -192 1230
rect -158 1196 -146 1230
rect -204 1190 -146 1196
rect -198 1158 -152 1190
rect -198 758 48 1158
rect 2 726 48 758
rect 2 680 102 726
rect 266 640 300 1271
rect 827 1230 885 1236
rect 827 1196 839 1230
rect 873 1196 885 1230
rect 827 1190 885 1196
rect 833 1158 879 1190
rect 361 758 371 1158
rect 423 758 433 1158
rect 619 758 629 1158
rect 681 758 879 1158
rect 266 606 414 640
rect -197 88 -1 488
rect 51 88 61 488
rect 247 88 257 488
rect 309 88 319 488
rect -198 87 47 88
rect -198 56 -152 87
rect -204 50 -146 56
rect -204 16 -192 50
rect -158 16 -146 50
rect -204 10 -146 16
rect 380 -25 414 606
rect 584 520 678 566
rect 632 488 678 520
rect 632 88 878 488
rect 832 56 878 88
rect 826 50 884 56
rect 826 16 838 50
rect 872 16 884 50
rect 826 10 884 16
rect 368 -31 426 -25
rect 368 -65 380 -31
rect 414 -65 426 -31
rect 368 -71 426 -65
<< via1 >>
rect 371 758 423 1158
rect 629 758 681 1158
rect -1 88 51 488
rect 257 88 309 488
<< metal2 >>
rect 371 1158 423 1168
rect 371 649 423 758
rect 627 1158 683 1168
rect 627 748 683 758
rect 257 597 423 649
rect -3 488 53 498
rect -3 78 53 88
rect 257 488 309 597
rect 257 78 309 88
<< via2 >>
rect 627 758 629 1158
rect 629 758 681 1158
rect 681 758 683 1158
rect -3 88 -1 488
rect -1 88 51 488
rect 51 88 53 488
<< metal3 >>
rect 617 1158 693 1163
rect 617 758 627 1158
rect 683 758 693 1158
rect 617 753 693 758
rect 625 655 685 753
rect -5 591 685 655
rect -5 493 55 591
rect -13 488 63 493
rect -13 88 -3 488
rect 53 88 63 488
rect -13 83 63 88
use sky130_fd_pr__nfet_01v8_8UMB6F  sky130_fd_pr__nfet_01v8_8UMB6F_0
timestamp 1729195750
transform 1 0 340 0 1 958
box -344 -288 344 288
use sky130_fd_pr__nfet_01v8_8UMB6F  sky130_fd_pr__nfet_01v8_8UMB6F_1
timestamp 1729195750
transform 1 0 340 0 1 288
box -344 -288 344 288
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_0
timestamp 1729189750
transform 1 0 -131 0 1 958
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_1
timestamp 1729189750
transform 1 0 812 0 1 958
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_2
timestamp 1729189750
transform 1 0 811 0 1 288
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_3
timestamp 1729189750
transform 1 0 -131 0 1 288
box -73 -226 73 226
<< labels >>
flabel metal2 396 711 396 711 0 FreeSans 320 0 0 0 RS
port 2 nsew
flabel metal1 25 703 25 703 0 FreeSans 320 0 0 0 D3
port 3 nsew
flabel metal3 655 625 655 625 0 FreeSans 320 0 0 0 D4
port 4 nsew
flabel metal1 281 1221 281 1221 0 FreeSans 320 0 0 0 GND
port 5 nsew
<< end >>
