magic
tech sky130A
magscale 1 2
timestamp 1729239979
<< nwell >>
rect -267 827 987 2045
<< nsubdiff >>
rect -231 1975 -171 2009
rect 891 1975 951 2009
rect -231 1953 -197 1975
rect 917 1953 951 1975
rect -231 897 -197 923
rect 917 897 951 923
rect -231 863 -171 897
rect 891 863 951 897
<< nsubdiffcont >>
rect -171 1975 891 2009
rect -231 923 -197 1953
rect 917 923 951 1953
rect -171 863 891 897
<< poly >>
rect -62 1863 30 1879
rect -62 1829 -46 1863
rect -12 1829 30 1863
rect -62 1813 30 1829
rect 0 1782 30 1813
rect 720 1863 812 1879
rect 720 1829 762 1863
rect 796 1829 812 1863
rect 720 1813 812 1829
rect 720 1782 750 1813
rect 0 1057 30 1088
rect -62 1041 30 1057
rect -62 1007 -46 1041
rect -12 1007 30 1041
rect -62 991 30 1007
rect 720 1057 750 1088
rect 720 1041 812 1057
rect 720 1007 762 1041
rect 796 1007 812 1041
rect 720 991 812 1007
<< polycont >>
rect -46 1829 -12 1863
rect 762 1829 796 1863
rect -46 1007 -12 1041
rect 762 1007 796 1041
<< locali >>
rect -231 1975 -171 2009
rect 891 1975 951 2009
rect -231 1953 -197 1975
rect 917 1953 951 1975
rect -62 1829 -46 1863
rect -12 1829 4 1863
rect 746 1829 762 1863
rect 796 1829 812 1863
rect -46 1782 -12 1829
rect 762 1780 796 1829
rect -46 1041 -12 1088
rect 762 1041 796 1088
rect -62 1007 -46 1041
rect -12 1007 4 1041
rect 746 1007 762 1041
rect 796 1007 812 1041
rect -231 897 -197 923
rect 917 897 951 923
rect -231 863 -171 897
rect 891 863 951 897
<< viali >>
rect 181 1975 533 2009
rect -46 1829 -12 1863
rect 762 1829 796 1863
rect -46 1007 -12 1041
rect 762 1007 796 1041
<< metal1 >>
rect 169 2009 545 2015
rect 169 1975 181 2009
rect 533 1975 545 2009
rect 169 1969 545 1975
rect -58 1863 0 1869
rect -58 1829 -46 1863
rect -12 1829 0 1863
rect -58 1823 0 1829
rect -46 1782 -12 1823
rect 99 1820 109 1872
rect 167 1820 177 1872
rect 257 1820 267 1872
rect 325 1820 335 1872
rect 415 1820 425 1872
rect 483 1820 493 1872
rect 573 1820 583 1872
rect 641 1820 651 1872
rect 750 1863 808 1869
rect 750 1829 762 1863
rect 796 1829 808 1863
rect 750 1823 808 1829
rect 762 1782 796 1823
rect -52 1770 82 1782
rect 668 1770 802 1782
rect -52 1594 33 1770
rect 85 1594 95 1770
rect -52 1582 82 1594
rect 94 1492 104 1544
rect 162 1492 172 1544
rect 200 1453 234 1770
rect 339 1594 349 1770
rect 401 1594 411 1770
rect 264 1495 274 1547
rect 330 1495 340 1547
rect 410 1495 420 1547
rect 476 1495 486 1547
rect 516 1453 550 1770
rect 655 1594 665 1770
rect 717 1594 802 1770
rect 668 1582 802 1594
rect 578 1492 588 1544
rect 646 1492 656 1544
rect 200 1425 550 1453
rect 94 1324 104 1380
rect 160 1324 170 1380
rect -52 1276 82 1288
rect -52 1100 33 1276
rect 85 1100 95 1276
rect 200 1100 234 1425
rect 262 1326 272 1378
rect 330 1326 340 1378
rect 410 1326 420 1378
rect 478 1326 488 1378
rect 339 1100 349 1276
rect 401 1100 411 1276
rect 516 1100 550 1425
rect 580 1326 590 1378
rect 646 1326 656 1378
rect 668 1276 802 1288
rect 655 1100 665 1276
rect 717 1100 802 1276
rect -52 1088 82 1100
rect 668 1088 802 1100
rect -46 1047 -12 1088
rect -58 1041 0 1047
rect -58 1007 -46 1041
rect -12 1007 0 1041
rect -58 1001 0 1007
rect 99 998 109 1050
rect 167 998 177 1050
rect 257 998 267 1050
rect 325 998 335 1050
rect 415 998 425 1050
rect 483 998 493 1050
rect 573 998 583 1050
rect 641 998 651 1050
rect 762 1047 796 1088
rect 750 1041 808 1047
rect 750 1007 762 1041
rect 796 1007 808 1041
rect 750 1001 808 1007
<< via1 >>
rect 109 1820 167 1872
rect 267 1820 325 1872
rect 425 1820 483 1872
rect 583 1820 641 1872
rect 33 1594 85 1770
rect 104 1492 162 1544
rect 349 1594 401 1770
rect 274 1495 330 1547
rect 420 1495 476 1547
rect 665 1594 717 1770
rect 588 1492 646 1544
rect 104 1324 160 1380
rect 33 1100 85 1276
rect 272 1326 330 1378
rect 420 1326 478 1378
rect 349 1100 401 1276
rect 590 1326 646 1378
rect 665 1100 717 1276
rect 109 998 167 1050
rect 267 998 325 1050
rect 425 998 483 1050
rect 583 998 641 1050
<< metal2 >>
rect -138 1918 392 1952
rect -138 960 -104 1918
rect 109 1872 167 1882
rect 109 1810 167 1820
rect 267 1872 325 1882
rect 267 1810 325 1820
rect 358 1780 392 1918
rect 425 1872 483 1882
rect 425 1810 483 1820
rect 583 1872 641 1882
rect 583 1810 641 1820
rect 31 1770 87 1780
rect 31 1584 87 1594
rect 349 1770 401 1780
rect 349 1584 401 1594
rect 663 1770 719 1780
rect 663 1584 719 1594
rect 104 1544 162 1554
rect 104 1456 162 1492
rect 274 1551 330 1561
rect 274 1485 330 1495
rect 420 1551 476 1561
rect 420 1485 476 1495
rect 588 1544 646 1554
rect 588 1456 646 1492
rect 104 1422 646 1456
rect 104 1380 160 1390
rect 104 1314 160 1324
rect 272 1378 330 1422
rect 272 1316 330 1326
rect 420 1378 478 1422
rect 420 1316 478 1326
rect 590 1378 646 1388
rect 590 1312 646 1322
rect 33 1276 85 1286
rect 33 1090 85 1100
rect 347 1276 403 1286
rect 347 1090 403 1100
rect 665 1276 717 1286
rect 665 1090 717 1100
rect 42 960 76 1090
rect 109 1050 167 1060
rect 109 988 167 998
rect 267 1050 325 1060
rect 267 988 325 998
rect 425 1050 483 1060
rect 425 988 483 998
rect 583 1050 641 1060
rect 583 988 641 998
rect 674 960 708 1090
rect -138 926 708 960
<< via2 >>
rect 31 1594 33 1770
rect 33 1594 85 1770
rect 85 1594 87 1770
rect 663 1594 665 1770
rect 665 1594 717 1770
rect 717 1594 719 1770
rect 274 1547 330 1551
rect 274 1495 330 1547
rect 420 1547 476 1551
rect 420 1495 476 1547
rect 104 1324 160 1380
rect 590 1326 646 1378
rect 590 1322 646 1326
rect 347 1100 349 1276
rect 349 1100 401 1276
rect 401 1100 403 1276
<< metal3 >>
rect 29 1898 890 1958
rect 29 1775 89 1898
rect 661 1775 721 1898
rect 21 1770 97 1775
rect 21 1594 31 1770
rect 87 1594 97 1770
rect 21 1589 97 1594
rect 653 1770 729 1775
rect 653 1594 663 1770
rect 719 1594 729 1770
rect 653 1589 729 1594
rect 262 1551 340 1556
rect 262 1495 274 1551
rect 330 1495 340 1551
rect 262 1467 340 1495
rect 410 1551 488 1556
rect 410 1495 420 1551
rect 476 1495 488 1551
rect 410 1467 488 1495
rect 94 1407 656 1467
rect 94 1380 172 1407
rect 94 1324 104 1380
rect 160 1324 172 1380
rect 94 1319 172 1324
rect 578 1378 656 1407
rect 578 1322 590 1378
rect 646 1322 656 1378
rect 578 1317 656 1322
rect 337 1276 413 1281
rect 337 1100 347 1276
rect 403 1100 413 1276
rect 337 1095 413 1100
rect 345 973 405 1095
rect 830 973 890 1898
rect 345 913 890 973
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729231575
transform 1 0 15 0 1 1188
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729231575
transform 1 0 735 0 1 1682
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729231575
transform 1 0 735 0 1 1188
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_6
timestamp 1729231575
transform 1 0 15 0 1 1682
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_VQXX7L  sky130_fd_pr__pfet_01v8_VQXX7L_0
timestamp 1729224175
transform 1 0 533 0 1 1188
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_VQXX7L  sky130_fd_pr__pfet_01v8_VQXX7L_1
timestamp 1729224175
transform 1 0 533 0 1 1682
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_VQXX7L  sky130_fd_pr__pfet_01v8_VQXX7L_6
timestamp 1729224175
transform 1 0 217 0 1 1188
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_VQXX7L  sky130_fd_pr__pfet_01v8_VQXX7L_7
timestamp 1729224175
transform 1 0 217 0 1 1682
box -223 -200 223 200
<< labels >>
flabel viali 347 1992 347 1992 0 FreeSans 320 0 0 0 VDD
port 3 nsew
flabel metal3 303 1472 303 1472 0 FreeSans 320 0 0 0 VIP
port 4 nsew
flabel metal2 454 1397 454 1397 0 FreeSans 320 0 0 0 VIN
port 5 nsew
flabel metal1 533 1556 533 1556 0 FreeSans 320 0 0 0 S
port 6 nsew
flabel metal2 -121 943 -121 943 0 FreeSans 320 0 0 0 OUT
port 12 nsew
flabel metal3 861 1929 861 1929 0 FreeSans 320 0 0 0 D6
port 14 nsew
<< end >>
