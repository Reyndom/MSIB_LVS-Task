magic
tech sky130A
magscale 1 2
timestamp 1729428971
<< viali >>
rect 395 1163 553 1197
rect 1186 1163 1344 1197
rect 1977 1163 2135 1197
rect 395 142 553 176
rect 1186 142 1344 176
rect 1977 142 2135 176
<< metal1 >>
rect 263 1197 2266 1233
rect 263 1163 395 1197
rect 553 1163 1186 1197
rect 1344 1163 1977 1197
rect 2135 1163 2266 1197
rect 263 1136 2266 1163
rect 376 639 386 691
rect 491 639 501 691
rect 562 645 1282 684
rect 1353 646 2073 685
rect 2134 638 2144 690
rect 2249 638 2259 690
rect 263 176 2266 203
rect 263 142 395 176
rect 553 142 1186 176
rect 1344 142 1977 176
rect 2135 142 2266 176
rect 263 106 2266 142
<< via1 >>
rect 386 639 491 691
rect 2144 638 2249 690
<< metal2 >>
rect 386 691 491 701
rect 2144 691 2249 700
rect 491 690 2249 691
rect 491 639 2144 690
rect 386 629 491 639
rect 2144 628 2249 638
use inverter  x1
timestamp 1729366069
transform 1 0 53 0 1 2350
box 210 -2244 632 -1117
use inverter  x2
timestamp 1729366069
transform 1 0 844 0 1 2350
box 210 -2244 632 -1117
use inverter  x3
timestamp 1729366069
transform 1 0 1635 0 1 2350
box 210 -2244 632 -1117
<< labels >>
flabel metal1 336 1179 336 1179 0 FreeSans 320 0 0 0 VDD
port 1 nsew
flabel metal1 335 153 335 153 0 FreeSans 320 0 0 0 GND
port 2 nsew
flabel via1 2197 663 2197 663 0 FreeSans 320 0 0 0 OUT
port 4 nsew
<< end >>
