magic
tech sky130A
magscale 1 2
timestamp 1729132732
<< error_p >>
rect -36 281 36 287
rect -36 247 -24 281
rect -36 241 36 247
rect -36 -247 36 -241
rect -36 -281 -24 -247
rect -36 -287 36 -281
<< nwell >>
rect -134 -300 134 300
<< pmos >>
rect -40 -200 40 200
<< pdiff >>
rect -98 188 -40 200
rect -98 -188 -86 188
rect -52 -188 -40 188
rect -98 -200 -40 -188
rect 40 188 98 200
rect 40 -188 52 188
rect 86 -188 98 188
rect 40 -200 98 -188
<< pdiffc >>
rect -86 -188 -52 188
rect 52 -188 86 188
<< poly >>
rect -40 281 40 297
rect -40 247 -24 281
rect 24 247 40 281
rect -40 200 40 247
rect -40 -247 40 -200
rect -40 -281 -24 -247
rect 24 -281 40 -247
rect -40 -297 40 -281
<< polycont >>
rect -24 247 24 281
rect -24 -281 24 -247
<< locali >>
rect -40 247 -24 281
rect 24 247 40 281
rect -86 188 -52 204
rect -86 -204 -52 -188
rect 52 188 86 204
rect 52 -204 86 -188
rect -40 -281 -24 -247
rect 24 -281 40 -247
<< viali >>
rect -24 247 24 281
rect -86 -188 -52 188
rect 52 -188 86 188
rect -24 -281 24 -247
<< metal1 >>
rect -36 281 36 287
rect -36 247 -24 281
rect 24 247 36 281
rect -36 241 36 247
rect -92 188 -46 200
rect -92 -188 -86 188
rect -52 -188 -46 188
rect -92 -200 -46 -188
rect 46 188 92 200
rect 46 -188 52 188
rect 86 -188 92 188
rect 46 -200 92 -188
rect -36 -247 36 -241
rect -36 -281 -24 -247
rect 24 -281 36 -247
rect -36 -287 36 -281
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.4 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
